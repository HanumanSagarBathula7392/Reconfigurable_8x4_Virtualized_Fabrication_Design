-- Company: 
-- Engineer: 
-- 
-- Create Date: 04/29/2024 01:06:19 PM
-- Design Name: 
-- Module Name: TOPMODULE_TB - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.NUMERIC_STD.ALL;
use ieee.std_logic_unsigned.all;
use std.env.finish;
use work.custom_pack.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity TOPMODULE_TB is
--  Port ( );
end TOPMODULE_TB;

architecture Behavioral of TOPMODULE_TB is
      constant dw: integer:=4;
      constant dws: integer:=5;
      constant dwm: integer:=2;
      constant rows: integer:=4;
      constant cols: integer:=4;
signal  A,B :  ARR_1D(0 to COLS-1) (DW-1 downto 0);
signal Y :  ARRAY_2D(0 to ROWS-1,0 to COLS-1) (DW-1 downto 0);
signal CLK:  std_logic:='0';
signal W_ENA,W_ENB,W_ENOP,W_ENY:  ARR_EN2D(0 to ROWS-1,0 to COLS-1);
signal SELMA,SELMB:  ARRAY_2D(0 to ROWS-1,0 to COLS-1)(DWM-1 downto 0);  
signal SELCU :  ARRAY_2D(0 to ROWS-1,0 to COLS-1)(DWS-1 downto 0);

begin

gm_i : entity work.TopModule

generic map(dw =>dw,dws=>dws,dwm=>dwm,rows=>rows,cols=>cols)
port map(A=>A,B=>B,Y=>Y,CLK=>CLK,
        W_ENA=>W_ENA,W_ENB=>W_ENB,W_ENY=>W_ENY,W_ENOP=>W_ENOP,
        SELMA=>SELMA,SELMB=>SELMB,SELCU=>SELCU);

CLK_PROC: process
begin
CLK<= not CLK after 5ns;
wait for 5 ns;
end process CLK_PROC;

stim:process
begin

---------------------RUN-1--------------------------
-------------EXTERNAL_INPUTS-------------------------
     A <= ("1010","1101","1010","1100");
     B <= ("0100","1011","1010","1010");
----------------------------------------------------
-----------------MUX_SELECTION--------------------
      SELMA <=(("00","01","01","00"),
                ("00","01","01","01"),
                ("00","10","10","01"),
                ("01","01","00","10"));
----------------------------------------------------
-------------------MUX_SELECTION--------------------               
      SELMB <=(("00","00","01","01"),
                ("00","00","00","01"),
                ("01","00","01","00"),
                ("00","10","01","00"));
------------------------------------------------------
------------------CU_SELECTION-----------------------                 
      SELCU <=(("00111","01000","00110","10011"),
                ("10010","10100","01110","01100"),
                ("00101","10101","00011","00001"),
                ("10011","01101","01000","00010"));
----------------------------------------------------
------------------ENABLE----------------------------
W_ENA <=(('0','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
W_ENB <=(('0','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
W_ENOP <=(('0','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
W_ENY <=(('0','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
 wait for 10 ns;
----------------------------------------------------
----------------------------------------------------
W_ENA <=(('1','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
W_ENB <=(('1','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('0','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
 wait for 20 ns;
----------------------------------------------------
----------------------------------------------------
W_ENA <=(('1','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
W_ENB <=(('1','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
 wait for 20 ns;
----------------------------------------------------
----------------------------------------------------
W_ENA <=(('1','1','1','1'),
        ('1','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
W_ENB <=(('1','1','1','1'),
        ('1','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
 wait for 20 ns;
----------------------------------------------------
W_ENA <=(('1','1','1','1'),
        ('1','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
W_ENB <=(('1','1','1','1'),
        ('1','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
 wait for 20 ns;
----------------------------------------------------
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'),
        ('0','0','0','0'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'),
        ('0','0','0','0'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','0','0','0'),
        ('0','0','0','0'),
        ('0','0','0','0'));
 wait for 20 ns; 
----------------------------------------------------
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'),
        ('0','0','0','0'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'),
        ('0','0','0','0'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'),
        ('0','0','0','0'));
 wait for 20 ns; 
---------------------------------------------------- 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'),
        ('0','0','0','0'));
 wait for 20 ns; 
---------------------------------------------------- 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'));
 wait for 20 ns; 
---------------------------------------------------- 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'));
 wait for 20 ns; 
---------------------------------------------------- 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
 wait for 20 ns; 
------------------------------------------------------ 
---------------------RUN-2--------------------------
-----------------MUX_SELECTION--------------------
      SELMA <=(("01","01","10","10"),
                ("00","01","01","01"),
                ("01","10","00","01"),
                ("00","00","00","01"));
----------------------------------------------------
-------------------MUX_SELECTION--------------------               
      SELMB <=(("01","10","01","01"),
                ("00","00","00","00"),
                ("00","00","01","00"),
                ("01","10","10","10"));
------------------------------------------------------
------------------CU_SELECTION-----------------------                 
      SELCU <=(("00100","00101","00011","01000"),
                ("00111","01100","00110","01110"),
                ("10010","01011","01000","00001"),
                ("01001","10101","10001","10100"));
                wait for 20 ns; 
----------------------------------------------------
------------------ENABLE----------------------------
W_ENA <=(('0','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENB <=(('0','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENOP <=(('0','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
 wait for 20 ns; 
------------------------------------------------------ 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('0','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
 wait for 20 ns; 
------------------------------------------------------ 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
 wait for 20 ns; 
------------------------------------------------------ 
W_ENA <=(('1','0','0','0'),
        ('0','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENB <=(('1','0','0','0'),
        ('0','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENOP <=(('1','0','0','0'),
        ('0','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
 wait for 20 ns; 
------------------------------------------------------ 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','0','0','0'),
        ('0','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
 wait for 20 ns; 
------------------------------------------------------ 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
 wait for 20 ns; 
------------------------------------------------------ 
W_ENA <=(('1','1','1','1'),
        ('1','0','0','0'),
        ('0','1','1','1'),
        ('1','1','1','1'));
W_ENB <=(('1','1','1','1'),
        ('1','0','0','0'),
        ('0','1','1','1'),
        ('1','1','1','1'));
W_ENOP <=(('1','1','1','1'),
        ('1','0','0','0'),
        ('0','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
 wait for 20 ns; 
------------------------------------------------------ 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','0','0','0'),
        ('0','1','1','1'),
        ('1','1','1','1'));
 wait for 20 ns; 
------------------------------------------------------ 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
 wait for 20 ns; 
------------------------------------------------------ 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'),
        ('0','1','1','1'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'),
        ('0','1','1','1'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'),
        ('0','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
 wait for 20 ns; 
------------------------------------------------------ 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'),
        ('0','1','1','1'));       
 wait for 20 ns; 
------------------------------------------------------ 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));      
 wait for 20 ns; 
------------------------------------------------------ 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));      
 wait for 20 ns; 
------------------------------------------------------ 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','0','0','0'));      
 wait for 20 ns; 
------------------------------------------------------ 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));      
 wait for 20 ns; 
------------------------------------------------------ 
W_ENA <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENB <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENOP <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));
W_ENY <=(('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'),
        ('1','1','1','1'));      
 wait for 20 ns; 
------------------------------------------------------ 
finish;    
 end process;
end Behavioral;
